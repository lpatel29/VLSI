module hello_world ;

initial begin
  $display ("Hello World by Linux");
  #10 $finish;
end

endmodule // End of Module hello_world
